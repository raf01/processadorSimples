module ULA (regA, regB, opcode, clock);

endmodule
