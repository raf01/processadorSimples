module UnidadeDeControle(opcode,rd,we);

input opcode;
output reg rd,we;
// fazer enable para o buffer de saida
always @(opcode)
begin
rd = 1'b0;
we = 1'b0;

	case(opcode)
		4'b0000:		//saida 0
			begin
				rd = 1'b0;
				we = 1'b0;
			end
		4'b0001:		//soma
			begin
				rd = 1'b0;
				we = 1'b0;

			end
		4'b0010:		//subtrai
			begin
				rd = 1'b0;
				we = 1'b0;
			end
		4'b0011:		//multiplica�ao
			begin
				rd = 1'b0;
				we = 1'b0;
			end
		4'b0100:		//divisao
			begin
				rd = 1'b0;
				we = 1'b0;
			end
		4'b0101:		//and
			begin
				rd = 1'b0;
				we = 1'b0;
			end
		4'b0110:		//or
			begin
				rd = 1'b0;
				we = 1'b0;
			end
		4'b0111:		//not
			begin
				rd = 1'b0;
				we = 1'b0;
			end
		4'b1000:		//xor
			begin
				rd = 1'b0;
				we = 1'b0;
			end
		4'b1001:		//xnor
			begin
				rd = 1'b0;		
				we = 1'b0;
			end
		4'b1010:		// Armazena o conteudo de a na saida da ULA
			begin
				rd = 1'b0;
				we = 1'b1; 
			end
		4'b1011:		// Armazena o conteudo de a na saida da ULA
			begin
				rd = 1'b0;
				we = 1'b1;
			end
		default:
			begin
				rd = 1'b0;
				we = 1'b0;
			
			end
	endcase
end 

endmodule 